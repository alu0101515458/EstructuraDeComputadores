module sum4(output wire[3:0] S, output wire c_out, input wire[3:0] A, input wire[3:0] B, input wire c_in)

  ul4 ul4_1();
  ul4 ul4_2();
  ul4 ul4_3();
  ul4 ul4_4();

endmodule